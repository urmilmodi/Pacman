`timescale 1ns / 1ns // `timescale time_unit/time_precision
module seg7_HEX0 (input [3:0]SW, output [6:0] HEX0);
    /*
        0  1  2  3  4  5  6
    0 - 0, 0, 0, 0, 0, 0, 1
    1 - 1, 0, 0, 1, 1, 1, 1
    2 - 0, 0, 1, 0, 0, 1, 0
    3 - 0, 0, 0, 0, 1, 1, 0
    4 - 1, 0, 0, 1, 1, 0, 0
    5 - 0, 1, 0, 0, 1, 0, 0
    6 - 0, 1, 0, 0, 0, 0, 0
    7 - 0, 0, 0, 1, 1, 1, 1
    8 - 0, 0, 0, 0, 0, 0, 0
    9 - 0, 0, 0, 1, 1, 0, 0
    A - 0, 0, 0, 1, 0, 0, 0
    b - 1, 1, 0, 0, 0, 0, 0
    C - 0, 1, 1, 0, 0, 0, 1
    d - 1, 0, 0, 0, 0, 1, 0
    E - 0, 1, 1, 0, 0, 0, 0
    F - 0, 1, 1, 1, 0, 0, 0
    */

    assign HEX0[0] = (~ SW[0] & ~ SW[1] & ~ SW[2] & SW[3]) | (~ SW[0] & SW[1] & ~ SW[2] & ~ SW[3]) | (SW[0] & ~ SW[1] & SW[2] & SW[3]) | (SW[0] & SW[1] & ~ SW[2] & SW[3]);
    assign HEX0[1] = (SW[0] & SW[1] & SW[2] & SW[3]) | (SW[0] & SW[1] & SW[2] & ~ SW[3]) | (SW[0] & SW[1] & ~ SW[2] & ~ SW[3]) | (SW[0] & ~ SW[1] & SW[2] & SW[3]) | (~ SW[0] & SW[1] & SW[2] & ~ SW[3]) | (~ SW[0] & SW[1] & ~ SW[2] & SW[3]);
    assign HEX0[2] = (SW[0] & SW[1] & SW[2] & SW[3]) | (SW[0] & SW[1] & SW[2] & ~ SW[3]) | (SW[0] & SW[1] & ~ SW[2] & ~ SW[3]) | (~ SW[0] & ~ SW[1] & SW[2] & ~ SW[3]);
    assign HEX0[3] = (SW[0] & SW[1] & SW[2] & SW[3]) | (SW[0] & ~ SW[1] & SW[2] & ~ SW[3]) | (SW[0] & ~ SW[1] & ~ SW[2] & SW[3]) | (~ SW[0] & SW[1] & SW[2] & SW[3]) | (~ SW[0] & SW[1] & ~ SW[2] & ~ SW[3]) | (~ SW[0] & ~ SW[1] & ~ SW[2] & SW[3]);
    assign HEX0[4] = (SW[0] & ~ SW[1] & ~ SW[2] & SW[3]) | (~ SW[0] & SW[1] & SW[2] & SW[3]) | (~ SW[0] & SW[1] & ~ SW[2] & SW[3]) | (~ SW[0] & SW[1] & ~ SW[2] & ~ SW[3]) | (~ SW[0] & ~ SW[1] & SW[2] & SW[3]) | (~ SW[0] & ~ SW[1] & ~ SW[2] & SW[3]);
    assign HEX0[5] = (SW[0] & SW[1] & ~ SW[2] & SW[3]) | (~ SW[0] & SW[1] & SW[2] & SW[3]) | (~ SW[0] & ~ SW[1] & SW[2] & SW[3]) | (~ SW[0] & ~ SW[1] & SW[2] & ~ SW[3]) | (~ SW[0] & ~ SW[1] & ~ SW[2] & SW[3]);
    assign HEX0[6] = (SW[0] & SW[1] & ~ SW[2] & ~ SW[3]) | (~ SW[0] & SW[1] & SW[2] & SW[3]) | (~ SW[0] & ~ SW[1] & ~ SW[2] & SW[3]) | (~ SW[0] & ~ SW[1] & ~ SW[2] & ~ SW[3]);
endmodule